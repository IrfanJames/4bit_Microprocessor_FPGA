module test_Cruncher();
	reg clk;
	wire Op_Code_Leds;
	
	initial
	begin
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
		clk = 0; #10;	clk = 1; #10;
	end
	
endmodule