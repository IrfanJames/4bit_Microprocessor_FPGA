//////////////////////////////////////////////////////////////////////////
// DFF for Cout of ALU

module D_ff (clk, in, out);
	input clk, in;
	output reg out;
	
	always @(posedge clk)
	begin
		if (clk)	out <= in;
	end
endmodule
//////////////////////////////////////////////////////////////////////////
